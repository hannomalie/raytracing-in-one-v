module main

struct World {
	sky Sky [required]
	objects []Hittable [required]
}

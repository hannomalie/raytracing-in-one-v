module main

fn degrees_to_radians(degrees f64) f64 {
	pi := 3.1415926535897932385
	return degrees * pi / 180.0
}
